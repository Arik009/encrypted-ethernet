`include "util.vh"
localparam BYTE_LEN = 8;

localparam PACKET_BUFFER_SIZE = 4096;
// taken from ip summary
localparam PACKET_BUFFER_READ_LATENCY = 2;

localparam PACKET_SYNTH_ROM_SIZE = 4096;
localparam PACKET_SYNTH_ROM_LATENCY = 2;

localparam SYNC_DELAY_LEN = 3;
