`include "util.vh"
localparam BYTE_LEN = 8;
localparam PACKET_BUFFER_SIZE = 4096;
// taken from ip summary
localparam PACKET_BUFFER_READ_LATENCY = 2;
